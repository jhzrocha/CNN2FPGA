
    LIBRARY ieee;
    USE ieee.std_logic_1164.ALL;

    PACKAGE types_pkg IS
type t_i_IN_DATA_poolingOperator_6_8_10 is array (0 to 5) of std_logic_vector(7 downto 0);

    END PACKAGE types_pkg;